* C:\Users\anjan\Desktop\Semester 4\Principles Of communication\PSPice\DSB.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 22 19:01:09 2021



** Analysis setup **
.tran 0ns 3m
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "DSB.net"
.INC "DSB.als"


.probe


.END
