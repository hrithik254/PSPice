* C:\Users\anjan\Desktop\Semester 4\Principles Of communication\PSPice\AM1.sch

* Schematics Version 9.1 - Web Update 1
* Sun Apr 04 23:05:12 2021



** Analysis setup **
.tran 0ns 1ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "AM1.net"
.INC "AM1.als"


.probe


.END
